library verilog;
use verilog.vl_types.all;
entity \SRA\ is
    port(
        x               : in     vl_logic_vector(31 downto 0);
        y               : in     vl_logic_vector(31 downto 0);
        \out\           : out    vl_logic_vector(31 downto 0)
    );
end \SRA\;
