library verilog;
use verilog.vl_types.all;
entity tlib_svh_unit is
end tlib_svh_unit;
