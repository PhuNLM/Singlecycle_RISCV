library verilog;
use verilog.vl_types.all;
entity singlecycle_vlg_vec_tst is
end singlecycle_vlg_vec_tst;
